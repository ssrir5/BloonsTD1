module life_counter(input logic )


endmodule