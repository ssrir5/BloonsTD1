module monkey_rom_backup( input [9:0] addressX, addressY,
								output data
								);
			
logic [4:0] X_bits, Y_bits;
logic [31:0] data_array;
			
assign X_bits = addressX[4:0];					 
assign Y_bits = addressY[4:0];				
	// ROM definition				
	logic [0:31][0:31] ROM = {
//         01234567890123456789012345678901
//                   1111111111222222222233
       32'b00000000000000011000000000000000, // 0 
       32'b00000000000111111111100000000000, // 1
       32'b00000000001111111111110000000000, // 2
       32'b00000000011111111111111000000000, // 3
       32'b00000000111111111111111100000000, // 4
       32'b00000001111111111111111110000000, // 5
       32'b00000011111111111111111111000000, // 6
       32'b00000111111111111111111111100000, // 7
       32'b00001111111111111111111111110000, // 8
       32'b00011111111111111111111111111000, // 9
       32'b00111111111111111111111111111100, // 10
       32'b01111111111111111111111111111110, // 11
       32'b11111111111111111111111111111111, // 12
       32'b11111111111111111111111111111111, // 13
       32'b11111111111111111111111111111111, // 14
       32'b01111111111111111111111111111110, // 15 
       32'b00011111111111111111111111111000, // 16
       32'b00000000000000000000000000000000, // 17
       32'b00000000000000000000000000000000, // 18
       32'b00000000000000000000000000000000, // 19
       32'b00000000000000000000000000000000, // 20
       32'b00000000000000000000000000000000, // 21
       32'b00000000000000000000000000000000, // 22
       32'b00000000000000000000000000000000, // 23
       32'b00000000000000000000000000000000, // 24
       32'b00000000000000000000000000000000, // 25
       32'b00000000000000000000000000000000, // 26
       32'b00000000000000000000000000000000, // 27
       32'b00000000000000000000000000000000, // 28
       32'b00000000000000000000000000000000, // 29
       32'b00000000000000000000000000000000, // 30
       32'b00000000000000000000000000000000, // 31
//         01234567890123456789012345678901
//                   1111111111222222222233
        };

	assign data_array = ROM[Y_bits];
	assign data = data_array[31-X_bits];
	

endmodule  